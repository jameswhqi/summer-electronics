// Tracking logic module
module Tracking
(
    
);

endmodule
module Pintest (
    input in,
    output reg out
);

    always @(*)
        out = in;

endmodule